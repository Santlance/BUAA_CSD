`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    10:52:52 11/08/2018 
// Design Name: 
// Module Name:    P1_11_1 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module P1_11_1(
		input clk,
		input clr,
		input [7:0] in,
		output reg out = 0
    );
	integer state = 0,bracket = 0;
	parameter  null = 0,

endmodule
