`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    10:43:42 10/07/2018 
// Design Name: 
// Module Name:    counter 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module counter(
    input clk,
    input rst_n,
    output [3:0] cnt 
    );
	 reg [3:0] count;
	 assign cnt=count;
	always@(posedge clk,negedge rst_n)
	begin 
	if(!rst_n)
	count<=0;
	else
	count<=count+1'b1;
	end

endmodule
