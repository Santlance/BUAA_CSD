`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    13:16:26 10/07/2018 
// Design Name: 
// Module Name:    sample 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////

//���Դ��ԵĽ�ģ�鹦�ܷ�Ϊ�������֣���������߼��ġ�����ʱ���߼��ġ��Լ�������ģ�������
//��������߼���ʹ��������ֵ���assign,assign���Ҳ��������������䣬ͨ������߼����ֶ�wire�ͱ�������������ֵ��Ҳ����ָ����ε����������������
//assign ��������һ��wire�ͱ������ұ���һ������߼��ı��ʽ��ͨ������߼��������ź�����������ٽ��õ��Ľ�������ұ�
//����������ݲ����������Ļ���ϵͳĬ����wire��
//verilog�е������������ͣ�wire �� reg
module sample(input clk);
	
	wire a;//��Ӧ��·ͼ�еĵ��ߣ�һ�������źţ�һ������źţ��������ܴ洢����
	reg b;//reg�ǼĴ������ͣ���Ӧ��·�еļĴ��������������д洢����
	//assign signal = expression;
	
	//ʱ���߼����֣�����ʱ���߼�������Ҫ���̿飬����initial��always��
	
	//initial����Ҫ�����ڳ���ʼʱ��ʼ�����������������������Ϊ��������ź�
	//ע�������begin end�ǿ�ı�־���൱��C�еĴ�����
	initial begin
	b = 0;
	end
	
	//always����Ҫ���ڷ�������в��ϼ������������������ʱ���Ὺʼִ�п��ڵĴ��룬����ʵ����ͨ���Ǽ���λ�仯
	//���б����ж������ʱ����������һ���������always�飬�����ָ��posedge��negede,�źŵ��κα仯���ᴥ�������д��@*���κα����ı仯���ᴥ��
	always @(posedge clk)begin
	b=~b;
	end
	//��һ��д��,�����ڱ仯��
	always #5 b=~b;//�����#5������ÿ���ʱ�䵥λ�󴥷�����
	
	
	//���һ��ģ������������ģ�飬����һ����·�л����������ӵ�·
	wire x,y,z;
	//Ҫָ��ģ����,�൱��һ�����ͣ�����һ���������ͺͱ�������Ȼ��Ҫ��ʵ����,ע�ⶥ��ģ�鲻���ٱ��ģ����ʵ����
	AndGate and1(x.y,z);//λ��ӳ��һһ��Ӧ
	AndGate and2(.b(x),.c(z));//��ӳ�䣬��.�����˿�֮������ӣ���ʱ����˳�����⣬��ʽΪ  .�˿������ź�����,�Ƽ�ʹ�ã�
	
	
endmodule
