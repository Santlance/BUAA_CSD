`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    20:24:09 10/29/2014 
// Design Name: 
// Module Name:    decoder 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module decoder(decoder_out,waddr,we);
		output[31:0] decoder_out;
		input[4:0] waddr;
		input we;
		reg [31:0] decoder_out;
		//input overflow;
		always @ (waddr or we)    
				//if ((we == 0) || (overflow == 1))
				if (we == 0)
						decoder_out = 32'h00000000;
				else
				case(waddr)
						5'd0:  decoder_out=32'b0000_0000_0000_0000_0000_0000_0000_0001;
						5'd1:  decoder_out=32'b0000_0000_0000_0000_0000_0000_0000_0010;
						5'd2:  decoder_out=32'b0000_0000_0000_0000_0000_0000_0000_0100;
						5'd3:  decoder_out=32'b0000_0000_0000_0000_0000_0000_0000_1000;
						5'd4:  decoder_out=32'b0000_0000_0000_0000_0000_0000_0001_0000;
						5'd5:  decoder_out=32'b0000_0000_0000_0000_0000_0000_0010_0000;
						5'd6:  decoder_out=32'b0000_0000_0000_0000_0000_0000_0100_0000;
						5'd7:  decoder_out=32'b0000_0000_0000_0000_0000_0000_1000_0000;
						5'd8:  decoder_out=32'b0000_0000_0000_0000_0000_0001_0000_0000;
						5'd9:  decoder_out=32'b0000_0000_0000_0000_0000_0010_0000_0000;
						5'd10: decoder_out=32'b0000_0000_0000_0000_0000_0100_0000_0000;
						5'd11: decoder_out=32'b0000_0000_0000_0000_0000_1000_0000_0000;
						5'd12: decoder_out=32'b0000_0000_0000_0000_0001_0000_0000_0000;
						5'd13: decoder_out=32'b0000_0000_0000_0000_0010_0000_0000_0000;
						5'd14: decoder_out=32'b0000_0000_0000_0000_0100_0000_0000_0000;
						5'd15: decoder_out=32'b0000_0000_0000_0000_1000_0000_0000_0000;
						5'd16: decoder_out=32'b0000_0000_0000_0001_0000_0000_0000_0000;
						5'd17: decoder_out=32'b0000_0000_0000_0010_0000_0000_0000_0000;
						5'd18: decoder_out=32'b0000_0000_0000_0100_0000_0000_0000_0000;
						5'd19: decoder_out=32'b0000_0000_0000_1000_0000_0000_0000_0000;
						5'd20: decoder_out=32'b0000_0000_0001_0000_0000_0000_0000_0000;
						5'd21: decoder_out=32'b0000_0000_0010_0000_0000_0000_0000_0000;
						5'd22: decoder_out=32'b0000_0000_0100_0000_0000_0000_0000_0000;
						5'd23: decoder_out=32'b0000_0000_1000_0000_0000_0000_0000_0000;
						5'd24: decoder_out=32'b0000_0001_0000_0000_0000_0000_0000_0000;
						5'd25: decoder_out=32'b0000_0010_0000_0000_0000_0000_0000_0000;
						5'd26: decoder_out=32'b0000_0100_0000_0000_0000_0000_0000_0000;
						5'd27: decoder_out=32'b0000_1000_0000_0000_0000_0000_0000_0000;
						5'd28: decoder_out=32'b0001_0000_0000_0000_0000_0000_0000_0000;
						5'd29: decoder_out=32'b0010_0000_0000_0000_0000_0000_0000_0000;
						5'd30: decoder_out=32'b0100_0000_0000_0000_0000_0000_0000_0000;
						5'd31: decoder_out=32'b1000_0000_0000_0000_0000_0000_0000_0000;
				endcase
endmodule