`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    23:48:46 10/21/2018 
// Design Name: 
// Module Name:    seven_digit 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module seven_digit(
	input x3,x2,x1,x0,
	output a,b,c,d,e,f,g
    );
	assign a=(!x3&&!x2&&!x1&&!x0)||(!x3&&!x2&&x1&&!x0)||(!x3&&!x2&&x1&&x0)||(!x3&&x2&&!x1&&x0)||(!x3&&x2&&x1&&!x0)||
	(!x3&&x2&&x1&&x0)||(x3&&!x2&&!x1&&!x0)||(x3&&!x2&&!x1&&x0)||(x3&&!x2&&x1&&!x0)||(x3&&x2&&!x1&&!x0)||(x3&&x2&&x1&&!x0)||
	(x3&&x2&&x1&&x0);
	
	assign b=(!x3&&!x2&&!x1&&!x0)||(!x3&&x2&&!x1&&!x0)||(!x3&&x2&&!x1&&x0)||(!x3&&x2&&x1&&!x0)||(x3&&!x2&&!x1&&!x0)||
	(x3&&!x2&&!x1&&x0)||(x3&&!x2&&x1&&!x0)||(x3&&!x2&&x1&&x0)||(x3&&x2&&!x1&&!x0)||(x3&&x2&&x1&&!x0)||(x3&&x2&&x1&&x0);
	
	assign c=(!x3&&!x2&&!x1&&!x0)||(!x3&&!x2&&x1&&!x0)||(!x3&&x2&&x1&&!x0)||(x3&&!x2&&!x1&&!x0)||(x3&&!x2&&x1&&!x0)||
	(x3&&!x2&&x1&&x0)||(x3&&x2&&!x1&&!x0)||(x3&&x2&&!x1&&x0)||(x3&&x2&&x1&&!x0)||(x3&&x2&&x1&&x0);
	
	assign d=(!x3&&!x2&&!x1&&!x0)||(!x3&&!x2&&x1&&!x0)||(!x3&&!x2&&x1&&x0)||(!x3&&x2&&!x1&&x0)||(!x3&&x2&&x1&&!x0)||
	(x3&&!x2&&!x1&&!x0)||(x3&&!x2&&!x1&&x0)||(x3&&!x2&&x1&&x0)||(x3&&x2&&!x1&&!x0)||(x3&&x2&&!x1&&x0)||(x3&&x2&&x1&&!x0);
	
	assign e=(!x3&&!x2&&!x1&&!x0)||(!x3&&!x2&&!x1&&x0)||(!x3&&!x2&&x1&&x0)||(!x3&&x2&&!x1&&!x0)||(!x3&&x2&&!x1&&x0)||
	(!x3&&x2&&x1&&!x0)||(!x3&&x2&&x1&&x0)||(x3&&!x2&&!x1&&!x0)||(x3&&!x2&&!x1&&x0)||(x3&&!x2&&x1&&!x0)||(x3&&!x2&&x1&&x0)||
	(x3&&x2&&!x1&&x0);
	
	assign f=(!x3&&!x2&&!x1&&!x0)||(!x3&&!x2&&!x1&&x0)||(!x3&&!x2&&x1&&!x0)||(!x3&&!x2&&x1&&x0)||(!x3&&x2&&!x1&&!x0)||
	(!x3&&x2&&x1&&x0)||(x3&&!x2&&!x1&&!x0)||(x3&&!x2&&!x1&&x0)||(x3&&!x2&&x1&&!x0)||(x3&&x2&&!x1&&x0);
	
	assign g=(!x3&&!x2&&x1&&!x0)||(!x3&&!x2&&x1&&x0)||(!x3&&x2&&!x1&&!x0)||(!x3&&x2&&!x1&&x0)||(!x3&&x2&&x1&&!x0)||
	(x3&&!x2&&!x1&&!x0)||(x3&&!x2&&!x1&&x0)||(x3&&!x2&&x1&&!x0)||(x3&&!x2&&x1&&x0)||(x3&&x2&&!x1&&x0)||(x3&&x2&&x1&&!x0)||
	(x3&&x2&&x1&&x0);

endmodule
