`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    12:49:51 11/25/2018 
// Design Name: 
// Module Name:    MUXALUIN 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module MUXALUIN(
	 input [31:0] out32,// 32
	 input [31:0] regdata2,// 32
	 input alusrc,// 1
	 
	 output [31:0] aluoprand_b// 32
    );


endmodule
