`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    12:49:40 11/25/2018 
// Design Name: 
// Module Name:    MUXREGIN 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module MUXREGIN(
	 input [4:0] rt,// 5
	 input [4:0] rd,// 5
	 input jal,// 1
	 input regdst,// 1
	 
	 output [4:0] regaddr// 5
    );


endmodule
